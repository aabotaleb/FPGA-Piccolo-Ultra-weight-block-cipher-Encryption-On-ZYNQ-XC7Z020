library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is
type ciphered_data is array (32 downto 0) of std_logic_vector(63 downto 0);
end constants;